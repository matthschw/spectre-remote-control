// Copied from CMOS Analog Circuit Design by Phillip E. Allen and Douglas R. Holberg
// Oxford University Press, Inc. , 2012
simulator lang=spice

.SUBCKT OPAMP 1 2 6 8 9
M1 4 2 3 3 NMOS1 W = 3U L = 1U AD = 18P AS = 18P PD = 18U PS =
+ 18U
M2 5 1 3 3 NMOS1 W = 3U L = 1U AD = 18P AS = 18P PD = 18U PS =
+ 18U
M3 4 4 8 8 PMOS1 W = 15U L = 1U AD = 90P AS = 90P PD = 42U PS = 42U
M4 5 4 8 8 PMOS1 W = 15U L = 1U AD = 90P AS = 90P PD = 42U PS = 42U
M5 3 7 9 9 NMOS1 W = 4.5U L = 1U AD = 27P AS = 27P PD = 21U PS = 21U
M6 6 5 8 8 PMOS1 W = 94U L = 1U AD = 564P AS = 564P PD = 200U PS = 200U
M7 6 7 9 9 NMOS1 W = 14U L = 1U AD = 84P AS = 84P PD = 40U PS = 40U
M8 7 7 9 9 NMOS1 W = 4.5U L = 1U AD = 27P AS = 27P PD = 21U PS = 21U
CC 5 6 3.0P
.MODEL NMOS1 NMOS VTO = 0.70 KP = 110U GAMMA = 0.4 LAMBDA = 0.04 PHI =
+ = 0.7 MJ = 0.5 MJSW = 0.38 CGBO = 700P CGSO = 220P CGDO = 220P CJ
+ = 770U CJSW = 380P LD = 0.016U TOX = 14N
.MODEL PMOS1 PMOS VTO = 20.7 KP = 50U GAMMA = 0.57 LAMBDA = 0.05 PHI
+ = 0.8 MJ = 0.5 MJSW = .35 CGBO = 700P CGSO = 220P CGDO = 220P CJ
+ = 560U CJSW = 350P LD = 0.014U TOX = 14N
IBIAS 8 7 30U
.ENDS

VIN1 1 0 DC 0 AC 1.0
VDD 4 0 DC 2.5
VSS 0 5 DC 2.5
VIN 2 2 0 DC 0
CL 3 0 10P
X1 1 2 3 4 5 OPAMP

.OP
.TF V(3) VIN1
.DC VIN1 20.005 0.005 100U
.AC DEC 10 1 10MEG
.END
